module mips_top
(input clk, rst, output [31:0] pc_current, instr, alu_out, wd_dm, rd_dm);
    wire we_dm;
    mips      MIPS (.clk(clk), .rst(rst), .instr(instr), .rd_dm(rd_dm), .we_dm(we_dm), .pc_current(pc_current), .alu_out(alu_out), .wd_dm(wd_dm));
    imem #(32)IMEM (.a(pc_current[7:2]), .y(instr));
    dmem #(32)DMEM (.clk(clk), .we(we_dm), .a(alu_out[5:0]), .d(wd_dm), .q(rd_dm));
endmodule

